`timescale 1ns / 1ps
`default_nettype none

module rasterize(
      input wire clk,
      input wire rst,
      input wire valid_in,
      input wire model_in,

      output logic valid,
      output logic pixel_out);




endmodule


`default_nettype wire
