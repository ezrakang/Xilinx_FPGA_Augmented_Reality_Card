`timescale 1ns / 1ps
`default_nettype none

module 3d_to_2d(
      input wire clk,
      input wire rst,
      input wire valid_in,
      input wire [63:0] model_in,
      input wire camera_loc,

      output logic valid,
      output logic model_out);




endmodule


`default_nettype wire
